-- Copyright (C) 2018  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.

-- Generated by Quartus Prime Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition
-- Created on Fri Oct 25 09:21:57 2024

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY maquina_estados00 IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        enable : IN STD_LOGIC := '0';
        sentido : IN STD_LOGIC := '0';
        saida1 : OUT STD_LOGIC;
        saida2 : OUT STD_LOGIC
    );
END maquina_estados00;

ARCHITECTURE BEHAVIOR OF maquina_estados00 IS
    TYPE type_fstate IS (s0,s1,s2,s3);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,enable,sentido)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= s0;
            saida1 <= '0';
            saida2 <= '0';
        ELSE
            saida1 <= '0';
            saida2 <= '0';
            CASE fstate IS
                WHEN s0 =>
                    IF (NOT((enable = '1'))) THEN
                        reg_fstate <= s0;
                    ELSIF (((enable = '1') AND (sentido = '1'))) THEN
                        reg_fstate <= s1;
                    ELSIF (((enable = '1') AND NOT((sentido = '1')))) THEN
                        reg_fstate <= s3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= s0;
                    END IF;

                    saida1 <= '1';

                    saida2 <= '1';
                WHEN s1 =>
                    IF (NOT((enable = '1'))) THEN
                        reg_fstate <= s1;
                    ELSIF (((enable = '1') AND (sentido = '1'))) THEN
                        reg_fstate <= s2;
                    ELSIF (((enable = '1') AND NOT((sentido = '1')))) THEN
                        reg_fstate <= s0;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= s1;
                    END IF;

                    saida1 <= '1';

                    saida2 <= '0';
                WHEN s2 =>
                    IF (NOT((enable = '1'))) THEN
                        reg_fstate <= s2;
                    ELSIF (((enable = '1') AND (sentido = '1'))) THEN
                        reg_fstate <= s3;
                    ELSIF (((enable = '1') AND NOT((sentido = '1')))) THEN
                        reg_fstate <= s1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= s2;
                    END IF;

                    saida1 <= '0';

                    saida2 <= '1';
                WHEN s3 =>
                    IF (NOT((enable = '1'))) THEN
                        reg_fstate <= s3;
                    ELSIF (((enable = '1') AND (sentido = '1'))) THEN
                        reg_fstate <= s0;
                    ELSIF (((enable = '1') AND NOT((sentido = '1')))) THEN
                        reg_fstate <= s2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= s3;
                    END IF;

                    saida1 <= '0';

                    saida2 <= '0';
                WHEN OTHERS => 
                    saida1 <= 'X';
                    saida2 <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
