-- Copyright (C) 2018  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.


-- Generated by Quartus Prime Version 18.1 (Build Build 625 09/12/2018)
-- Created on Fri Nov 01 09:24:13 2024

robo_seguidor_linha_exemplo robo_seguidor_linha_exemplo_inst
(
	.reset(reset_sig) ,	// input  reset_sig
	.clock(clock_sig) ,	// input  clock_sig
	.sensord(sensord_sig) ,	// input  sensord_sig
	.sensore(sensore_sig) ,	// input  sensore_sig
	.ligamotordir(ligamotordir_sig) ,	// output  ligamotordir_sig
	.ligamotoresq(ligamotoresq_sig) ,	// output  ligamotoresq_sig
	.velmotordir(velmotordir_sig) ,	// output  velmotordir_sig
	.velmotoresq(velmotoresq_sig) 	// output  velmotoresq_sig
);

