-- Copyright (C) 2018  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.

-- Generated by Quartus Prime Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition
-- Created on Thu Oct 31 23:46:10 2024

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY atividade02_seguidor_linha IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        ligado : IN STD_LOGIC := '0';
        esgotou : IN STD_LOGIC := '0';
        sensor_esq : IN STD_LOGIC := '0';
        sensor_dir : IN STD_LOGIC := '0';
        motor_dir_full : OUT STD_LOGIC;
        motor_dir_half : OUT STD_LOGIC;
        motor_esq_full : OUT STD_LOGIC;
        motor_esq_half : OUT STD_LOGIC
    );
END atividade02_seguidor_linha;

ARCHITECTURE BEHAVIOR OF atividade02_seguidor_linha IS
    TYPE type_fstate IS (parado,frente,dir_half,esq_half,dir_full,esq_full);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,ligado,esgotou,sensor_esq,sensor_dir)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= parado;
            motor_dir_full <= '0';
            motor_dir_half <= '0';
            motor_esq_full <= '0';
            motor_esq_half <= '0';
        ELSE
            motor_dir_full <= '0';
            motor_dir_half <= '0';
            motor_esq_full <= '0';
            motor_esq_half <= '0';
            CASE fstate IS
                WHEN parado =>
                    IF ((NOT((sensor_dir = '1')) AND NOT((sensor_esq = '1')))) THEN
                        reg_fstate <= parado;
                    ELSIF ((((ligado = '1') AND (sensor_dir = '1')) AND (sensor_esq = '1'))) THEN
                        reg_fstate <= frente;
                    ELSIF ((((ligado = '1') AND NOT((sensor_dir = '1'))) AND (sensor_esq = '1'))) THEN
                        reg_fstate <= dir_full;
                    ELSIF ((((ligado = '1') AND (sensor_dir = '1')) AND NOT((sensor_esq = '1')))) THEN
                        reg_fstate <= esq_full;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= parado;
                    END IF;

                    motor_dir_half <= '0';

                    motor_dir_full <= '0';

                    motor_esq_full <= '0';

                    motor_esq_half <= '0';
                WHEN frente =>
                    IF ((((ligado = '1') AND NOT((sensor_dir = '1'))) AND (sensor_esq = '1'))) THEN
                        reg_fstate <= dir_full;
                    ELSIF ((((ligado = '1') AND (sensor_dir = '1')) AND NOT((sensor_esq = '1')))) THEN
                        reg_fstate <= esq_full;
                    ELSIF ((((ligado = '1') AND (sensor_dir = '1')) AND (sensor_esq = '1'))) THEN
                        reg_fstate <= frente;
                    ELSIF ((((ligado = '1') AND NOT((sensor_dir = '1'))) AND NOT((sensor_esq = '1')))) THEN
                        reg_fstate <= parado;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= frente;
                    END IF;

                    motor_dir_half <= '0';

                    motor_dir_full <= '1';

                    motor_esq_full <= '1';

                    motor_esq_half <= '0';
                WHEN dir_half =>
                    IF (((((ligado = '1') AND (esgotou = '1')) AND NOT((sensor_dir = '1'))) AND NOT((sensor_esq = '1')))) THEN
                        reg_fstate <= parado;
                    ELSIF (((((ligado = '1') AND NOT((esgotou = '1'))) AND (sensor_dir = '1')) AND (sensor_esq = '1'))) THEN
                        reg_fstate <= frente;
                    ELSIF (((((ligado = '1') AND NOT((esgotou = '1'))) AND NOT((sensor_dir = '1'))) AND NOT((sensor_esq = '1')))) THEN
                        reg_fstate <= dir_half;
                    ELSIF (((((ligado = '1') AND NOT((esgotou = '1'))) AND NOT((sensor_dir = '1'))) AND (sensor_esq = '1'))) THEN
                        reg_fstate <= dir_full;
                    ELSIF (((((ligado = '1') AND NOT((esgotou = '1'))) AND (sensor_dir = '1')) AND NOT((sensor_esq = '1')))) THEN
                        reg_fstate <= esq_full;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= dir_half;
                    END IF;

                    motor_dir_half <= '1';

                    motor_dir_full <= '0';

                    motor_esq_full <= '0';

                    motor_esq_half <= '0';
                WHEN esq_half =>
                    IF (((((ligado = '1') AND (esgotou = '1')) AND NOT((sensor_dir = '1'))) AND NOT((sensor_esq = '1')))) THEN
                        reg_fstate <= parado;
                    ELSIF (((((ligado = '1') AND NOT((esgotou = '1'))) AND (sensor_dir = '1')) AND (sensor_esq = '1'))) THEN
                        reg_fstate <= frente;
                    ELSIF (((((ligado = '1') AND NOT((esgotou = '1'))) AND NOT((sensor_dir = '1'))) AND NOT((sensor_esq = '1')))) THEN
                        reg_fstate <= esq_half;
                    ELSIF (((((ligado = '1') AND NOT((esgotou = '1'))) AND NOT((sensor_dir = '1'))) AND (sensor_esq = '1'))) THEN
                        reg_fstate <= dir_full;
                    ELSIF (((((ligado = '1') AND NOT((esgotou = '1'))) AND (sensor_dir = '1')) AND NOT((sensor_esq = '1')))) THEN
                        reg_fstate <= esq_full;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= esq_half;
                    END IF;

                    motor_dir_half <= '0';

                    motor_dir_full <= '0';

                    motor_esq_full <= '0';

                    motor_esq_half <= '1';
                WHEN dir_full =>
                    IF ((((ligado = '1') AND NOT((sensor_dir = '1'))) AND NOT((sensor_esq = '1')))) THEN
                        reg_fstate <= dir_half;
                    ELSIF ((((ligado = '1') AND (sensor_dir = '1')) AND (sensor_esq = '1'))) THEN
                        reg_fstate <= frente;
                    ELSIF ((((ligado = '1') AND NOT((sensor_dir = '1'))) AND (sensor_esq = '1'))) THEN
                        reg_fstate <= dir_full;
                    ELSIF ((((ligado = '1') AND (sensor_dir = '1')) AND NOT((sensor_esq = '1')))) THEN
                        reg_fstate <= esq_full;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= dir_full;
                    END IF;

                    motor_dir_half <= '0';

                    motor_dir_full <= '1';

                    motor_esq_full <= '0';

                    motor_esq_half <= '0';
                WHEN esq_full =>
                    IF ((((ligado = '1') AND NOT((sensor_dir = '1'))) AND NOT((sensor_esq = '1')))) THEN
                        reg_fstate <= esq_half;
                    ELSIF ((((ligado = '1') AND (sensor_dir = '1')) AND (sensor_esq = '1'))) THEN
                        reg_fstate <= frente;
                    ELSIF ((((ligado = '1') AND (sensor_dir = '1')) AND NOT((sensor_esq = '1')))) THEN
                        reg_fstate <= esq_full;
                    ELSIF ((((ligado = '1') AND NOT((sensor_dir = '1'))) AND (sensor_esq = '1'))) THEN
                        reg_fstate <= dir_full;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= esq_full;
                    END IF;

                    motor_dir_half <= '0';

                    motor_dir_full <= '0';

                    motor_esq_full <= '1';

                    motor_esq_half <= '0';
                WHEN OTHERS => 
                    motor_dir_full <= 'X';
                    motor_dir_half <= 'X';
                    motor_esq_full <= 'X';
                    motor_esq_half <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
