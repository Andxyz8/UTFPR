comparador_inst : comparador PORT MAP (
		dataa	 => dataa_sig,
		aeb	 => aeb_sig
	);
