-- megafunction wizard: %LPM_COUNTER%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: LPM_COUNTER 

-- ============================================================
-- File Name: divisor_barra.vhd
-- Megafunction Name(s):
-- 			LPM_COUNTER
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 18.1.0 Build 625 09/12/2018 SJ Lite Edition
-- ************************************************************


--Copyright (C) 2018  Intel Corporation. All rights reserved.
--Your use of Intel Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Intel Program License 
--Subscription Agreement, the Intel Quartus Prime License Agreement,
--the Intel FPGA IP License Agreement, or other applicable license
--agreement, including, without limitation, that your use is for
--the sole purpose of programming logic devices manufactured by
--Intel and sold by Intel or its authorized distributors.  Please
--refer to the applicable agreement for further details.


LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

LIBRARY lpm;
USE lpm.ALL;

ENTITY clock_barra IS
	PORT
	(
		clock		: IN STD_LOGIC ;
		q		: OUT STD_LOGIC_VECTOR (24 DOWNTO 0)
	);
END clock_barra;


ARCHITECTURE sincronizar OF clock_barra IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (24 DOWNTO 0);


	COMPONENT lpm_counter
		GENERIC (
			lpm_direction: STRING;
			lpm_port_updown: STRING;
			lpm_type: STRING;
			lpm_width: NATURAL
		);

		PORT (
			clock	: IN STD_LOGIC ;
			q	: OUT STD_LOGIC_VECTOR (24 DOWNTO 0)
		);
	END COMPONENT;


	BEGIN
		q <= sub_wire0(24 DOWNTO 0);

		LPM_COUNTER_component : LPM_COUNTER

		GENERIC MAP (
			lpm_direction => "UP",
			lpm_port_updown => "PORT_UNUSED",
			lpm_type => "LPM_COUNTER",
			lpm_width => 25
		)

		PORT MAP (
			clock => clock,
			q => sub_wire0
		);

END sincronizar;
