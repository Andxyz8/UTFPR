-- Copyright (C) 2018  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.


-- Generated by Quartus Prime Version 18.1 (Build Build 625 09/12/2018)
-- Created on Thu Oct 31 23:46:14 2024

atividade02_seguidor_linha atividade02_seguidor_linha_inst
(
	.reset(reset_sig) ,	// input  reset_sig
	.clock(clock_sig) ,	// input  clock_sig
	.ligado(ligado_sig) ,	// input  ligado_sig
	.esgotou(esgotou_sig) ,	// input  esgotou_sig
	.sensor_esq(sensor_esq_sig) ,	// input  sensor_esq_sig
	.sensor_dir(sensor_dir_sig) ,	// input  sensor_dir_sig
	.motor_dir_full(motor_dir_full_sig) ,	// output  motor_dir_full_sig
	.motor_dir_half(motor_dir_half_sig) ,	// output  motor_dir_half_sig
	.motor_esq_full(motor_esq_full_sig) ,	// output  motor_esq_full_sig
	.motor_esq_half(motor_esq_half_sig) 	// output  motor_esq_half_sig
);

