cont2_inst : cont2 PORT MAP (
		clock	 => clock_sig,
		q	 => q_sig
	);
