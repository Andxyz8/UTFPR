contador1_inst : contador1 PORT MAP (
		clock	 => clock_sig,
		q	 => q_sig
	);
