-- Copyright (C) 2018  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.

-- Generated by Quartus Prime Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition
-- Created on Fri Nov 01 09:18:36 2024

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY robo_seguidor_linha_exemplo IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        sensord : IN STD_LOGIC := '0';
        sensore : IN STD_LOGIC := '0';
        ligamotordir : OUT STD_LOGIC;
        ligamotoresq : OUT STD_LOGIC;
        velmotordir : OUT STD_LOGIC;
        velmotoresq : OUT STD_LOGIC
    );
END robo_seguidor_linha_exemplo;

ARCHITECTURE BEHAVIOR OF robo_seguidor_linha_exemplo IS
    TYPE type_fstate IS (nalinha,saidaesq,saidadir,foradalinha);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,sensord,sensore)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= nalinha;
            ligamotordir <= '0';
            ligamotoresq <= '0';
            velmotordir <= '0';
            velmotoresq <= '0';
        ELSE
            ligamotordir <= '0';
            ligamotoresq <= '0';
            velmotordir <= '0';
            velmotoresq <= '0';
            CASE fstate IS
                WHEN nalinha =>
                    IF (((sensord = '1') AND (sensore = '1'))) THEN
                        reg_fstate <= nalinha;
                    ELSIF (((sensord = '1') AND NOT((sensore = '1')))) THEN
                        reg_fstate <= saidaesq;
                    ELSIF ((NOT((sensord = '1')) AND (sensore = '1'))) THEN
                        reg_fstate <= saidadir;
                    ELSIF ((NOT((sensord = '1')) AND NOT((sensore = '1')))) THEN
                        reg_fstate <= foradalinha;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= nalinha;
                    END IF;

                    ligamotoresq <= '1';

                    ligamotordir <= '1';

                    velmotordir <= '1';

                    velmotoresq <= '1';
                WHEN saidaesq =>
                    IF (((sensord = '1') AND (sensore = '1'))) THEN
                        reg_fstate <= nalinha;
                    ELSIF ((NOT((sensord = '1')) AND NOT((sensore = '1')))) THEN
                        reg_fstate <= foradalinha;
                    ELSIF (((sensord = '1') AND NOT((sensore = '1')))) THEN
                        reg_fstate <= saidaesq;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= saidaesq;
                    END IF;

                    ligamotoresq <= '1';

                    ligamotordir <= '0';

                    velmotoresq <= '0';
                WHEN saidadir =>
                    IF (((sensord = '1') AND (sensore = '1'))) THEN
                        reg_fstate <= nalinha;
                    ELSIF ((NOT((sensord = '1')) AND NOT((sensore = '1')))) THEN
                        reg_fstate <= foradalinha;
                    ELSIF ((NOT((sensord = '1')) AND (sensore = '1'))) THEN
                        reg_fstate <= saidadir;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= saidadir;
                    END IF;

                    ligamotoresq <= '0';

                    ligamotordir <= '1';

                    velmotordir <= '0';
                WHEN foradalinha =>
                    IF ((NOT((sensord = '1')) AND NOT((sensore = '1')))) THEN
                        reg_fstate <= foradalinha;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= foradalinha;
                    END IF;

                    ligamotoresq <= '0';

                    ligamotordir <= '0';
                WHEN OTHERS => 
                    ligamotordir <= 'X';
                    ligamotoresq <= 'X';
                    velmotordir <= 'X';
                    velmotoresq <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
